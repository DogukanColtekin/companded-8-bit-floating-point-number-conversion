library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity elevenbittobcd is
    Port ( mult : in STD_LOGIC_VECTOR(10 downto 0);
           bcdbits : out STD_LOGIC_VECTOR(15 downto 0));
end elevenbittobcd;

architecture dataflow of elevenbittobcd is

begin

with mult select
    bcdbits <=
        "0000000000000000" when "00000000000",  
        "0000000000000001" when "00000000001",  
        "0000000000000010" when "00000000010",  
        "0000000000000011" when "00000000011",  
        "0000000000000100" when "00000000100",  
        "0000000000000101" when "00000000101",  
        "0000000000000110" when "00000000110",  
        "0000000000000111" when "00000000111",  
        "0000000000001000" when "00000001000",  
        "0000000000001001" when "00000001001",  
        "0000000000010000" when "00000001010",  
        "0000000000010001" when "00000001011",  
        "0000000000010010" when "00000001100",  
        "0000000000010011" when "00000001101",  
        "0000000000010100" when "00000001110", 
        "0000000000010101" when "00000001111",  
        "0000000000010110" when "00000010000",  
        "0000000000011000" when "00000010010",  
        "0000000000100000" when "00000010100",  
        "0000000000100010" when "00000010110",  
        "0000000000100100" when "00000011000",  
        "0000000000100110" when "00000011010",  
        "0000000000101000" when "00000011100",  
        "0000000000110000" when "00000011110",  
        "0000000000110010" when "00000100000", 
        "0000000000110110" when "00000100100",  
        "0000000001000000" when "00000101000",  
        "0000000001000100" when "00000101100",  
        "0000000001001000" when "00000110000",  
        "0000000001010010" when "00000110100", 
        "0000000001010110" when "00000111000",
        "0000000001100000" when "00000111100",  
        "0000000001100100" when "00001000000", 
        "0000000001110010" when "00001001000",
        "0000000010000000" when "00001010000",  
        "0000000010001000" when "00001011000",  
        "0000000010010110" when "00001100000",  
        "0000000100000100" when "00001101000", 
        "0000000100010010" when "00001110000",  
        "0000000100100000" when "00001111000",  
        "0000000100101000" when "00010000000",  
        "0000000101000100" when "00010010000",  
        "0000000101100000" when "00010100000",  
        "0000000101110110" when "00010110000",  
        "0000000110010010" when "00011000000", 
        "0000001000001000" when "00011010000", 
        "0000001000100100" when "00011100000",  
        "0000001001000000" when "00011110000", 
        "0000001001010110" when "00100000000",  
        "0000001010001000" when "00100100000",  
        "0000001100100000" when "00101000000",  
        "0000001101010010" when "00101100000", 
        "0000001110000100" when "00110000000", 
        "0000010000010110" when "00110100000", 
        "0000010001001000" when "00111000000",  
        "0000010010000000" when "00111100000",  
        "0000010100010010" when "01000000000", 
        "0000010101110110" when "01001000000",  
        "0000011001000000" when "01010000000",  
        "0000011100000100" when "01011000000",  
        "0000011101101000" when "01100000000",  
        "0000100000110010" when "01101000000",  
        "0000100010010110" when "01110000000",  
        "0000100101100000" when "01111000000",  
        "0001000000100100" when "10000000000",  
        "0001000101010010" when "10010000000",  
        "0001001010000000" when "10100000000",  
        "0001010000001000" when "10110000000",  
        "0001010100110110" when "11000000000",  
        "0001011001100100" when "11010000000",  
        "0001011110010010" when "11100000000", 
        "0001100100100000" when "11110000000", 
        "0000000000000000" when others;

end dataflow;